`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:51:06 06/18/2017 
// Design Name: 
// Module Name:    DECODE 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DECODE(
    output [31:0] instruction_in,
    output [31:0] data1_out,
    output [31:0] data2_out,
    output [5:0] opcode_out,
    output [5:0] funcode_out,
    input clock
    );


endmodule
